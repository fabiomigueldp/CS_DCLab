library ieee;use ieee.std_logic_1164.all;use ieee.numeric_std.all;entity jankenpon is port(A,B,C,D,H:in std_logic;HEX4:out std_logic_vector(6 downto 0));end;architecture a of jankenpon is constant L:std_logic_vector(223 downto 0):=x"00000000103CA4009207901E5240FFFFFFFFFFFFFFFFFFFFFFFFFFFF";begin HEX4<=L((to_integer(unsigned(H&A&B&C&D))*7+6)downto(to_integer(unsigned(H&A&B&C&D))*7));end;